.PARAM
+ LM1 = 7.6105e-07
+ LM2 = 5.9433e-07
+ LM3 = 1.1792e-06
+ WM1 = 8.0403e-05
+ WM2 = 4.2798e-05
+ WM3 = 9.1221e-06
+ Ib = 7.5191e-05
