.PARAM
+ LM1 = 7.7221e-07
+ LM2 = 6.4897e-07
+ LM3 = 1.1857e-06
+ WM1 = 8.0581e-05
+ WM2 = 3.9573e-05
+ WM3 = 8.1485e-06
+ Ib = 7.4531e-05
