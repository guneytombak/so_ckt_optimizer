.PARAM
+ LM1 = 3.5634e-07
+ LM2 = 6.871e-07
+ LM3 = 1.1732e-06
+ WM1 = 8.0447e-05
+ WM2 = 4.0685e-05
+ WM3 = 1.1646e-05
+ Ib = 7.525e-05
