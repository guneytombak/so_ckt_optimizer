.PARAM
+ LM1 = 7.2585e-07
+ LM2 = 6.9683e-07
+ LM3 = 1.1576e-06
+ WM1 = 7.9749e-05
+ WM2 = 4.0313e-05
+ WM3 = 4.6546e-06
+ Ib = 7.8837e-05
